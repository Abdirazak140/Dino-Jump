module HexDisplay();